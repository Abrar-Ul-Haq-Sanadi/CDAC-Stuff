library verilog;
use verilog.vl_types.all;
entity abc is
end abc;
