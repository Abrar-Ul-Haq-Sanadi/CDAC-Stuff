`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 18.05.2024 21:52:17
// Design Name: 
// Module Name: lab66_tb_101_Non_Overlap_OneHot_Encode_Moore
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module lab66_tb_101_Non_Overlap_OneHot_Encode_Moore(

    );
endmodule
