// DSCH3
// 10-07-2024 20:02:33
// C:\Users\vlsi\Desktop\CMOS\DSCH\Abu_Hash_schematic\inverter_sym.sch

module inverter_sym( clk1,out1);
 input clk1;
 output out1;
 wire ;
 not inv_1(out1,clk1);
endmodule
