// DSCH3
// 11-07-2024 19:31:03
// C:\Users\vlsi\Desktop\CMOS\DSCH\Abu_Hash_schematic\OR_Gate\or2_sym.sch

module or2_sym( in1,in2,out1);
 input in1,in2;
 output out1;
 wire ;
 or or2_1(out1,in1,in2);
endmodule
