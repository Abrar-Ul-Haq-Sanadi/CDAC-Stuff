CIRCUIT example
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
VA 9 0 PULSE(0.00 1.20 1.98N 0.02N 0.03N 1.97N 4.00N)
VB 11 0 PULSE(0.00 1.20 0.98N 0.03N 0.02N 0.98N 2.00N)
*
* List of nodes
* " xor2_Sum" corresponds to n�3
* "N4" corresponds to n�4
* "N5" corresponds to n�5
* " and2_Carry" corresponds to n�7
* "N8" corresponds to n�8
* "A" corresponds to n�9
* "B" corresponds to n�11
*
* MOS devices
MN1 0 4 3 0 N1  W= 0.24U L= 0.12U
MN2 9 11 4 0 N1  W= 0.24U L= 0.12U
MN3 0 9 5 0 N1  W= 0.24U L= 0.12U
MN4 0 8 7 0 N1  W= 0.24U L= 0.12U
MN5 10 9 8 0 N1  W= 0.24U L= 0.12U
MN6 0 11 10 0 N1  W= 0.24U L= 0.12U
MP1 1 4 3 1 P1  W= 0.72U L= 0.12U
MP2 5 11 4 1 P1  W= 0.72U L= 0.12U
MP3 1 9 5 1 P1  W= 0.72U L= 0.12U
MP4 1 8 7 1 P1  W= 0.72U L= 0.12U
MP5 8 9 1 1 P1  W= 0.72U L= 0.12U
MP6 1 11 8 1 P1  W= 0.72U L= 0.12U
*
C2 1 0  4.677fF
C3 3 0  0.819fF
C4 4 0  0.680fF
C5 5 0  0.524fF
C7 7 0  0.688fF
C8 8 0  0.706fF
C9 9 0  0.997fF
C10 10 0  0.090fF
C11 11 0  0.827fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.1N 5.00N
* (Pspice)
.PROBE
.END
