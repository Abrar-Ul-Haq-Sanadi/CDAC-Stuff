library verilog;
use verilog.vl_types.all;
entity phases_uvm_sv_unit is
end phases_uvm_sv_unit;
