CIRCUIT C:\Users\vlsi\Desktop\CMOS\DSCH\Abu_Hash_schematic\Cmos_lab_exam\exnor_layout.MSK
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
V~B 9 0 PULSE(0.00 1.20 0.48N 0.03N 0.03N 0.48N 1.00N)
VA 10 0 PULSE(0.00 1.20 0.23N 0.03N 0.03N 0.23N 0.50N)
V~A 11 0 PULSE(1.20 0.00 0.23N 0.03N 0.03N 0.23N 0.50N)
VB 12 0 PULSE(1.20 0.00 0.48N 0.03N 0.03N 0.48N 1.00N)
*
* List of nodes
* "Out" corresponds to n�3
* "N4" corresponds to n�4
* "N6" corresponds to n�6
* "N7" corresponds to n�7
* "~B" corresponds to n�9
* "A" corresponds to n�10
* "~A" corresponds to n�11
* "B" corresponds to n�12
*
* MOS devices
MN1 3 10 6 0 N1  W= 0.60U L= 0.12U
MN2 7 11 3 0 N1  W= 0.60U L= 0.12U
MN3 0 12 7 0 N1  W= 0.60U L= 0.12U
MN4 6 9 0 0 N1  W= 0.60U L= 0.12U
MP1 4 10 3 1 P1  W= 0.60U L= 0.12U
MP2 1 11 4 1 P1  W= 0.60U L= 0.12U
MP3 4 12 1 1 P1  W= 0.60U L= 0.12U
MP4 3 9 4 1 P1  W= 0.60U L= 0.12U
*
C2 1 0  0.950fF
C3 3 0  0.740fF
C4 4 0  0.480fF
C5 1 0  0.201fF
C6 6 0  0.493fF
C7 7 0  0.212fF
C9 9 0  0.132fF
C10 10 0  0.132fF
C11 11 0  0.132fF
C12 12 0  0.132fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.1N 5.00N
* (Pspice)
.PROBE
.END
