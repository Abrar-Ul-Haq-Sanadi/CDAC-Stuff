// Interface.sv
interface full_subtractor_if();
    logic a;
    logic b;
    logic bin;
    logic diff;
    logic bout;
endinterface