// DSCH3
// 07-08-2014 02:19:43 PM
// D:\installed program\DSCH\System\examples\flashMemory.sch

module flashMemory( );
 wire w2,w3,w4,w5,w6,w7,w8,w9;
 wire w10,w11,w12,w13,w14,w15;
//Warning: dgmos (dgmos) ignored 
//Warning: dgmos (dgmos) ignored 
//Warning: dgmos (dgmos) ignored 
//Warning: IO (Source) ignored 
//Warning: dgmos (dgmos) ignored 
//Warning: IO (Source) ignored 
//Warning: dgmos (dgmos) ignored 
//Warning: dgmos (dgmos) ignored 
//Warning: IO (0V) ignored 
//Warning: IO (HVDD) ignored 
//Warning: IO (0V) ignored 
//Warning: dgmos (dgmos) ignored 
//Warning: dgmos (dgmos) ignored 
//Warning: dgmos (dgmos) ignored 
endmodule

// Simulation parameters in Verilog Format

// Simulation parameters
