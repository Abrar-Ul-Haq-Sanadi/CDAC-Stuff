library verilog;
use verilog.vl_types.all;
entity adder_top_sv_unit is
end adder_top_sv_unit;
