library verilog;
use verilog.vl_types.all;
entity Uvm_phases_sv_unit is
end Uvm_phases_sv_unit;
