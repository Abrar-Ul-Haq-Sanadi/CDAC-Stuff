// DSCH3
// 11-07-2024 20:54:16
// C:\Users\vlsi\Desktop\CMOS\DSCH\Abu_Hash_schematic\AND_GATE\and2_symb.sch

module and2_symb( in1,in2,out1);
 input in1,in2;
 output out1;
 wire ;
 and and2_1(out1,in2,in1);
endmodule
