CIRCUIT example
*
* IC Technology: CMOS 0.12�m - 6 Metal
*
VDD 1 0 DC 1.20
*
* List of nodes
* "xor" corresponds to n�3
* "nxor" corresponds to n�4
* "N5" corresponds to n�5
* "inv" corresponds to n�7
* "a" corresponds to n�8
* "in" corresponds to n�9
* "b" corresponds to n�10
*
* MOS devices
MN1 0 4 3 0 N1  W= 0.24U L= 0.12U
MN2 8 10 4 0 N1  W= 0.24U L= 0.12U
MN3 0 8 5 0 N1  W= 0.24U L= 0.12U
MN4 0 9 7 0 N1  W= 0.24U L= 0.12U
MP1 1 4 3 1 P1  W= 0.72U L= 0.12U
MP2 5 10 4 1 P1  W= 0.72U L= 0.12U
MP3 1 8 5 1 P1  W= 0.72U L= 0.12U
MP4 1 9 7 1 P1  W= 0.72U L= 0.12U
*
C2 1 0  3.401fF
C3 3 0  0.524fF
C4 4 0  0.680fF
C5 5 0  0.524fF
C7 7 0  0.524fF
C8 8 0  0.480fF
C9 9 0  0.314fF
C10 10 0  0.314fF
*
* n-MOS Model 3 :
* low leakage
.MODEL N1 NMOS LEVEL=3 VTO=0.40 UO=600.000 TOX= 2.0E-9
+LD =0.000U THETA=0.500 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=120.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* p-MOS Model 3:
* low leakage
.MODEL P1 PMOS LEVEL=3 VTO=-0.45 UO=200.000 TOX= 2.0E-9
+LD =0.000U THETA=0.300 GAMMA=0.400
+PHI=0.200 KAPPA=0.060 VMAX=110.00K
+CGSO=100.0p CGDO=100.0p
+CGBO= 60.0p CJSW=240.0p
*
* Transient analysis
*
.TEMP 27.0
.TRAN 0.1N 5.00N
* (Pspice)
.PROBE
.END
